// TODO: revisar si es necesario el output de address
// error en address, definir otro nombre para el output 

module topRam(input logic clk, rst,
				  input logic [2:0] btn,
				  output [31:0] q,
				  output [15:0] address);
				  
logic wren;
logic [31:0] data;

ram mem(address, clk, data, wren, q);

write_mem escribir(btn, wren, address, data);


endmodule

module Testbench;
  //RandomNumberGenerator rng;

  initial begin
    // Simular durante un período de tiempo
    #1000;
    $finish;
  end
endmodule
